
`define max(a,b)((a) > (b) ? (a) : (b))
`define min(a,b)((a) < (b) ? (a) : (b))

module soc_rom
  #(parameter VECTOR_LENGTH = 'd512,
    parameter WORD_WIDTH = 'd16, // 8, 16 or 32
    parameter ADDR_WIDTH = ceil_log2(VECTOR_LENGTH))
   (
    output [WORD_WIDTH-1:0] data_o,
    input                   clk_i,
    input                   sel_i,
    input                   read_i,
    input [ADDR_WIDTH-1:0]  addr_i
    );

   function integer ceil_log2;
      input [31:0] arg;
      integer      i;
      begin
         ceil_log2 = 0;
         for (i = 0; i < 32; i = i + 1) begin
            if (arg > (1 << i))
              ceil_log2 = ceil_log2 + 1;
         end
      end
   endfunction

   wire [31:0] rdata32;
   wire [7:0]  addr;

   generate
      if (WORD_WIDTH == 'd8) begin : u_8bit
         reg byte_addr_q;

         assign data_o = byte_addr_q ? rdata32[15:8] : rdata32[7:0];
         assign addr = addr_i[`min(8,ADDR_WIDTH-1):1];

         always @(posedge clk_i) begin
            if (sel_i & read_i)
              byte_addr_q <= addr_i[0];
         end
      end else if (WORD_WIDTH == 'd16) begin : u_16bit
         assign data_o = rdata32[15:0];
         assign addr = addr_i[`min(7,ADDR_WIDTH-1):0];
      end else begin : u_32bit
         assign data_o = rdata32;
         assign addr = addr_i[`min(7,ADDR_WIDTH-1):0];
      end
   endgenerate

   localparam ROM_WORDS = (WORD_WIDTH == 'd32) ? 2 : 1;
   localparam ROM_BLOCKS = (((WORD_WIDTH == 'd8) ? (VECTOR_LENGTH+1)/2 : VECTOR_LENGTH)+255)/256;
   wire [16*ROM_BLOCKS*ROM_WORDS-1:0] rdata;
   wire [`max(ceil_log2(ROM_BLOCKS)-1, 0):0] block_addr;

   generate
      if (ROM_BLOCKS > 1) begin : u_multi_bank
         reg [ceil_log2(ROM_BLOCKS)-1:0] block_addr_q;

         assign block_addr = addr_i[ADDR_WIDTH-1 -:ceil_log2(ROM_BLOCKS)];
         assign rdata32[15:0] = rdata[16*ROM_WORDS*block_addr_q +:16];
         if (ROM_WORDS > 1) begin : u_high_word
            assign rdata32[31:16] = rdata[16*(ROM_WORDS*block_addr_q+1) +:16];
         end

         always @(posedge clk_i) begin
            if (sel_i & read_i)
              block_addr_q <= block_addr;
         end
      end else begin : u_single_bank
         assign block_addr = 0;
         assign rdata32[15:0] = rdata[15:0];
         if (ROM_WORDS > 1) begin : u_high_word
            assign rdata32[31:16] = rdata[31:16];
         end
      end
   endgenerate

   localparam [256*16*16-1:0] ROM_DATA = {256'hF879D288DA537D24E5B2B5F3E7B9291CB94FD333F808530DFB98D8E196DE6F3E,
                                          256'hDBE1B8E7CBC80A5436AEB5E3EAB52BC6730CC248434EBC8D71374DCF5762AEF3,
                                          256'h36DB27ADC1C169383F7F42DCFED1DF47113D72F5D0138332A69DADD90782F165,
                                          256'h1FD85FC0B91997EB62042641D64A897B524860AA9D0E6A1E536F2CC658D32323,
                                          256'h583031F1B2F42B6BA93DE369C7622FB8C19E14322D4C4224DCF4A19DFF9D4E32,
                                          256'h10A7C57A43E225F2E830B3718A1466D75300649B7C236ED8FB70304653CB6A2B,
                                          256'hC4BA12197D62FC029CB5499E717BD8876B793A8C17850FC6981D5253BC6EC86C,
                                          256'h25FC92D668F691C9E9860E7B91FD6CEBE9642998F0665ADB8F637CC0F5D95823,
                                          256'h2919156FA186F16D64AE1A42DB7CD26491E2C89764A57B5A7153C2387FEC3B32,
                                          256'hF114DB9289D14B1E5053EE1C2A9E1FE50A3085B50F4395A18B6FB4D4CF565FFD,
                                          256'h76619E87AF3102E1B30BE05C786D47ADCE47CFF8D7EE276D4A73DAC43BF50979,
                                          256'hDE61D4184EB76B59BF0D77E82C7AC9159EF82A48081B5804E994BFC280E0368B,
                                          256'h64590BFCD9F59E387C75672AEB618A1B9368475814CB1C07416DFF9A65E645E2,
                                          256'hAD6DCE3FB091BF91E527966A238CCD481CA9840AFF90FC111D80DDC624CB9016,
                                          256'h696AD1FAEC27A8D111E04C29C11B271B98DD34E52071E085FE0DE0619F796035,
                                          256'h35DCB6254B8EB75391FE0D578FC49AEECDE7E9EFEDE3C95C5D4097A8A9EDD0CB,
                                          256'h6494A012B5B84A961342C1E374CE8C0C9EDC89581A58E8C791D6C953F4A6E6FC,
                                          256'h9C62C41E53FD6F53A4D702801E6A588DBCAFB3978E71C9665A925FD3BB52EE6F,
                                          256'h699CE08667C639D1D63B05A43743175FD79C9250D22F8AD6726CC7F48AADD537,
                                          256'hA2F417AB5885B0D2D482415EB22AAAF3ED28656673F20CCA3DECDADDC12F9FC9,
                                          256'h7126334077B2D709299B429102A80948146E502FAE7E2E48A172D8E068AF1156,
                                          256'hE61303E6257993A00974466184169A59625CEF985B1858D746B867DF5D6F8AC9,
                                          256'hC67F0A01C2F9BD49C2809DF0FFE8D6C72CA9050FA05395916D718B182CFF5B44,
                                          256'h3705DC8F3EB4CC0A778054E5879642330BCA734F3758FB749C397E6EAE6C1A57,
                                          256'h4CE293504666BED1877FF1786220D7051CFCA554B94E983CF2BA47F4E8F54347,
                                          256'hBBADDE784A48D6952948FBB5B95F7FE7B7E32F3150A622FBDB26DC7083081C92,
                                          256'h53FF66A860B7616B3E17337925C686F1003687926504932290AB29FE4184D708,
                                          256'h949EA62C67D5012B198C08C97255A37DD48F972345B4A4D0348B5BFE9F0511C4,
                                          256'hB971B1FDF7F2AE716A4CFF5B9ADD1767DC7C9112DC4CCA429EF34D00DF6CBF4D,
                                          256'hDBFA79AF78EC322E813AB8500E46C76AA21868FDD19EF7E6BB1B5D82945C04C6,
                                          256'h7733A2F3AC6F7D5940173B316AD0F329EE309D3760F61174D46D3FFD8005B630,
                                          256'h8DD2BE7AE2140A5277658EACF0E59A7B2CA6530B098218DAC380F4DD3F0E7C10,
                                          256'hF84B074E8F774425A47C2F6C2D87D5110C1CE60E65871B7D75996D4C7EF73F6C,
                                          256'h7375289AD5881A471E134F1328DC6AA7D8FA83F5A836D3975F94C008F3BB5A93,
                                          256'hEEA4E68569925B59EE1FEF7D9DBA452B8CD93315B76F7312DA7A9CD44ED05CEB,
                                          256'hB51EDC25F9D40062859971146DE71D6063684AC03D00D2CBAF7AFE48BE9ECD57,
                                          256'hC51025C08EBC32B4B4A14C750946FAF02578FCD75B2776A8E9D6DF7159B917E5,
                                          256'h8438C92C37BCD4A944C2B6BE078197664CC9708F81B6A60B29A30EB8DDDF9929,
                                          256'hF7F52C824A6D4AD39884DD3842BAE49FF12ADDBFFD7B0AEF5E5119EEDDD8EB24,
                                          256'hE94F8EC5644B9F68A4F2C73654D6CC8A0D03E9FE7E96B388D773FF68E1F723B5,
                                          256'hBB7C2EF81F1375D74F8DCFA04E85572DE240D6BB1825F8083C8C4A53FC44FE8E,
                                          256'h1D3F7EC21D30D3EA0171421DE53BBCB3A31D5DD887D4230052499E86A8E22C92,
                                          256'hCFEFE1FE4C6C79015F2AF91778A946052989E83D74A0992CC50E52479DDBA61D,
                                          256'h210BD88CA2B72AC98E444B01FDBE021B38A041A9A1DDF9B3839D2F4D555C71E2,
                                          256'h7813AE88FD740DC58354AD8D986DF0716E7D1CF07F11EC773265C09ADBC4B86F,
                                          256'hFE5EA7DF4BB00130BA2DF27E0CF409C323CA3BB9FE65E733696618B56BF9B739,
                                          256'hE096710FBAA0E4526F5A4D55A0FA2A02A0759B3B3649F0526E11AC58A82102C2,
                                          256'h6581A9B3457EBB77C91225974A76F83EB5758912B6BBFA2CE4496E2B8445A157,
                                          256'hE28B70631F26FF6DA7AAFA5D5FB880207CFB2248EE93E13CAC1BF7F11C14EA5B,
                                          256'hC9D636524502D38685816CF46C04688411C2EF4E6B931F1F819F598000183ED6,
                                          256'hC1F4F04A3C4F6A17D77F0EA7CD6D63FD3E7B8FF5E2D1D9A374CC8F9BCDC47C0E,
                                          256'hFAE7601CA507378F618C0B5AFC6026179241B119E253A101D74AB9B266011BA0,
                                          256'hD7C69900DA93E4FC83077DE7C06C7805587A5F99C0440A9AC47626DC81F23EC3,
                                          256'h22AD6A901D6B5AB0A2CF3966EA2E0E6B9423AA968102AD29799D11A129C58913,
                                          256'h3186247853EB294AF7199B0C3C49C84EE6EAD14BDD4B8F3F4B8E0CC957B123C5,
                                          256'h16F3FF6710538F903A871CB3FDA5F701E46B94BD90C2F7043DD1BF9927AB72D2,
                                          256'h9BAFE3A9A2CAA4029A93134851BEB8C40D3C8ADACA8C374129DFABED897B685E,
                                          256'h5B42057595C81C457CF9F3E5BB70673C9AC852B38D0C4C291D1DCDF1EFFC5C06,
                                          256'h2F3161E0C220BD1B2DC051EB11FFAC36A05A086F15F6CA5BDB8E8346E93DFEA4,
                                          256'h66FCC276EEE8E8634761F084B3D26BBC6A96B2E2DFFB2657E16DF2973F0B1C52,
                                          256'hA05A44D19BD8F2D82E98C1A67F7C2E089188F091D740AA507C240E540E193E6D,
                                          256'h234042C6278063EC52DF8676E31B5F4C244514909B1B8239DFCF5F31D9BBE79E,
                                          256'h75F3289C1518C558051CB7DA6B1EFAB2D3D6B58886696C87247C5048C9E97318,
                                          256'h98AD95F03D7E94AA2FFE87D7AD7EDFB40881892B2E865556607878591F0AC591,
                                          256'h8DD182885C3C5557F7CE67B653C87D102D3F0586D09B41A3F74149B6348CE40A,
                                          256'h9BD229562BD029528ECA38E95A7C302062E30CB50A7CE9CF2AD8C1FF80DE04B3,
                                          256'h05C727E7AD4D2954DA098B8C2737B2D78E9DC5C51AAABB3B4508C6E1E1D5CB55,
                                          256'h7E22273FA02788002FCCD380ACA8335781FE131B2068805047DCF1158838C9A0,
                                          256'hD480C0D8C0F60A51A45C61A835B57E0E8C7E32827CE98A45326332FAD6F1BC5C,
                                          256'hFE0B6FB41EEB5B7719C5320F1A8841C83D67E36EED2991F1FDD7C61EF1A9790B,
                                          256'h15DEB8C7A800D80A54130E4A3AD6E86B461A038109B2DC60B5B412E448184D0B,
                                          256'h376A4ABE721C5EE40691F1DF3A226A048E25E1A638A6CCFE2CFB47278E82EE17,
                                          256'hF33E621B81ACF625BDFE7F135C80E17E54C2E5D6339EF75E49F67AB838DD332B,
                                          256'h027CAB476D7A04E4DC68377459D71260250D7D93ADC25B592DB40816E88F2ACC,
                                          256'h9C9C74B9E8FE9747089ECEB6EA0B084EB1A0C5D7CB8EB6401C5A81B4A918E43B,
                                          256'hD457CFB9D35D096E3E518C8359F9C935D658B6689B21EE7AA4C5118E496B6030,
                                          256'h374D4A45DC1C3E1273DCA47E5967232F339673BEA852DCAB28489647F26B5326,
                                          256'hFE635819200EC692126F21D283302D3CC79F63457CF889B08EB6DD2285E232A6,
                                          256'h4720DD7F5DC5BE4ACE402B9A0E4A4B1DFE70B5563A83B52FDB4C85794202404B,
                                          256'h3ED46367FE12C5B2A1D8A48CB970D1227B4892FF203DA7BBBBA7B6266F40AF03,
                                          256'h3682381DC1F5BD72267329526CD2C5292AA8F4121954A1B9361835AA5800822C,
                                          256'h33EC2F3A798D3C1BAF52E52FAD9275A6B345DD5C00F5C8D9BE181FD22C0C9099,
                                          256'hA67D4CECA602ECDFDB4789E34D3DBE6D705BD83A032B225530CBB21E4C76C0DA,
                                          256'h478A0A0202A49427BAFCBB2779AC058BF0040F4990BF5B7FA01D33173E200D4E,
                                          256'hAE3F772107AE018D48424753A5655E716921D40F32371E43506B4BA84D4F0871,
                                          256'h5E0A4CCC6C74CC5CE3C1A9FF9F26DB7CA7C836A3F225E2E40EF854BCDA190179,
                                          256'h00D684D2887A6CF1BA5E6EC976ABB7180653A1D8F46A753DC27B91854B4AF92F,
                                          256'h29BA1393A3AFAF2BCEF7EE9F05996BF1B99DD742FA44A6F29EA10D354FBBF20E,
                                          256'h3495D4B6F1E6CD252EBA826D97DF2DE732EDD73F41C70D6318364B58A049FAFA,
                                          256'h6A29EC823F2A3E31EB1CB822FC4B41E80641A8978C6FB912AFDD768630EC9D33,
                                          256'h85355ECA53795965373E63B34C8C6E0210E4CB1BDE1A43599DF7672A311B18CF,
                                          256'h5718149AF6EAD1833EEB773363323A2CCDAA451CCD23C5E7951BD3DB8D95175E,
                                          256'hAC9A3604F5DEEDB35D72CD6E962233052EF4468A3EA100FE1D969977F543F42C,
                                          256'h0B40602EB4FEFD0E55923E3CBDB22069C65E4AB4F66032E0CD5A148C3832C03D,
                                          256'h93B752F1C6F0B18D3647EAD1AF155AD78439AAF9BF3FC8889D556FDC8D55A472,
                                          256'hFE75448CFBC3040568154F51F9660F2CA2A3F68B06F7EBB3DF744C10A5A74A87,
                                          256'h7AFFEA8DAB2E6FD243AFBD5DAC0A21345BF3FB72D1346FE7AF9CEE2E488F57A4,
                                          256'h744488115DC16FC99ED2F24B8C4DD49118D2F555CB9F2E9E64F530B1CA51B84C,
                                          256'hE9F1F0F802E1EC588A80EAA80DBD90AE9ACDA0BBB65D0DB3191464ECEAFC2D40,
                                          256'hD731E40D607A68006391B76A58AB4D0FFBFFF0AFAFBCFA88DFEC081D197BB2EF,
                                          256'h41B814A61435BCEBA965F27EE21B822A768F20F1B1ABB85C3F66766DB5690755,
                                          256'h699D534F46ECF7343F87642932927B763B38B6F86336DB1A495FA8301DF14540,
                                          256'h50AB2B58FDE1E3E77C2F37C10651251C1ACFC5D051D61F7075ECB8B66FBB5D31,
                                          256'h12DE1A96D2F71F73D10D4A54DD6A0F6B233673B1050E8D48940E44A25EC29643,
                                          256'h278B3DDE9D56E3863AAFB3C2E20BD011543201B3EF52DCF6C046F83A8245F4CA,
                                          256'h02A7C66EC976F2E0982793CB670C2E91DF709D199C94F25BFABF891BAA288474,
                                          256'hD8B7155D225D9A89A520C8B7EA4690E4A4011DE84019DB9873DC11371D180C76,
                                          256'h535651698395FF154389F28849A17F6F505D13B3549B6032144143A30D50B3B9,
                                          256'h6A9A5A5511A4079886B359CB65590CD18A62154B1B44A32F83150683F31645A7,
                                          256'hFA43FE04D0E5F7487796AAB2CE234FF2F16C08B0F9F2C5F196AF6FAA04C6701D,
                                          256'hF6AFDD0D40C758EEADF1A3E777B11B56CD004C6B8FA3955FA9E3A61BA8F71859,
                                          256'h8EF95C8C8AA3F0CF49FD31B718D672AEC560F6FE32FF5E97C1BB3E016CC97870,
                                          256'hE0313CDEB1B743E4254778615A85D92B9295C54ED5DA6CF3A551A79A6BDB39D8,
                                          256'h693B2B49728D93EAC5033A49CEA34646E7A14D8DC0CAA4FEF05D387DF307A25C,
                                          256'hE50C675090E79F716B1C677269959D5473D46CAED5AD4FB371BF4C2AEF55228C,
                                          256'hF74FFDB9BFD8D3B17FA91E673E7B409B0BB196FC46071F07917454A3B0B45C85,
                                          256'h1ECB85730C06B34758739AAA8A8AC837F0CF68D6D1808140D8F62C6FD73911C6,
                                          256'h8703324C0AE98EEF77BE1072932A66622ED1D8942651ECCD4E0C875A85EBE9E5,
                                          256'hB34340D6CBEC8611C89FDC8421C34E5ED731203B5528429834759F69A9ED1FC0,
                                          256'h25B7E6C451F67EBB81EEA5E7085C1221958457E95BB1EDD5244C44B99FF33565,
                                          256'h7808BDE557B372A119FE75E35F25FB8332B23C14FF4408BCFD5F62376367ADFD,
                                          256'h5B9F5352EEE2DF688D1205583758692EA090B74C71E7D7657ED818BA7178CD9F,
                                          256'h0461FB33396266C9B4680BC884F4EF5E77CC0969BA3491AB4D2C852BAD979FB4,
                                          256'hB8339CF28D5357ECCC1D68BD1EE4A61EF3BF1A4DA2420E2F14E568B6FD5CE4EF,
                                          256'hC8F33BCEBA38E6D8ACA32A20AAA96EA454F7EB602228DD2AA3837A12DF82C4DE,
                                          256'h7727E8B872C2F0ABC173EC20A412F547393D2001A5C2C0835B253C107DD96E30,
                                          256'h6E37386B2EDFECEBDD7A3FC77FF3119A63B2225AAF96647487C1DC10BF8BB2E7,
                                          256'h502C44E16A96CC178EB542F680B6465A437F77D0FE9713E906D585F52B884EEB,
                                          256'h9BB5A2D0C5C14552149CE296C568E66FBC332A2A803D34EB4B4534B7CD8E50A7,
                                          256'hA1ED2F9A2281F22AEB54F388C043975EBC56B0710DC2EF40B14FC169AA57A5F5,
                                          256'h49BF753DD441C5417FE26AA8CBE353D4E1A319B1A3B801288B66E46C4155185A,
                                          256'hAC44BC4F0F73420FB0EEE150BFC418D7EEDED145CB2671AE752250F351AC5DF2,
                                          256'h985E739F09A971D216E3F115FD5A936C3F2B3A0156B0E8428775FC944E55CD8B,
                                          256'hB3C0A45F35A2E9F77739DA45B40576CE77D8133163B49487C992D694E8B17A2C,
                                          256'h020245CF12972585972BBEE75BD92C648A533DCCAC0799293819E72A92E1EB1F,
                                          256'h6B8726152847B3DFE6FC02C5AB66242BE27F529056081381042ADF0FDD3D5150,
                                          256'h499FB2669AD8C016BA4C9AA00F57352F2919B0472EC74CED74FE84686C467A66,
                                          256'h21F508B029C16A9862AFDDA518DC1D57F003C7FF273D9F2468CA8A54FC0AFCBF,
                                          256'h441C8E22EDB8E9D1B0E8957D1A6FE77C0BB28F6F8CCD5218B7D89FF9EB4B8E8C,
                                          256'h5CA9D233E18F414E02373C56BDBA34BE5ADE99C08A333941FBE97C79CAFC59DB,
                                          256'h56400934CAE27A9E20FCB50FD95D901830F0349B4FBD97FF11BF44DCDC1AC195,
                                          256'h51A41066C6520733490ED75A2092F1AA4895A1A7E9C217072DCD888FE950859D,
                                          256'h80B360454C5B61A5C0F692880EADED5F6B7F303E4C6D65BFD24CBDAF71EED3DF,
                                          256'hEF226E391B324FC8D26D0C255458A872DB1EAF974A33E4F0D5E46F3C9C8F3CB1,
                                          256'h0AC21D194128E54A0415CD1C6A0AF0C1B5A4C5D6C11D218AA223615FC9661DAB,
                                          256'hB2FCD2718339C4516812059638235CFEBAC3F1FB0BF1D26C84E15EF8FF33D7B6,
                                          256'hEBAA24502EDBD662C1118AE2DDEC61B299082A8567EA7D44A853A0F7DD71C25F,
                                          256'h81743003984812E9B445E2FBE97F2D164F04E987CA2CC77A858646AD16171F17,
                                          256'hD50392396598A5A82615A5FB633BDC34D993F0C31B3FFA43E4CE373B800DE378,
                                          256'hCAF2CE5BEDE6E2B51EF18582F5BE91543936D4C79F02C9FE10EF135F5856AE84,
                                          256'h271273C968AF080D63898A9931512F9AD9D924FECB6AA3502C54955F520D87A0,
                                          256'h755F430EE50D8840C274B1660E8B52107F73215FEF16318DF13160725A755724,
                                          256'hC17C69CF3C2838C1507E51700190136542A4B165F313BCDAF9677C686674D425,
                                          256'h7A2934CC8605F365F7D3F2D242C11ADCCB065C9CFDD2159B75CA253B5308F289,
                                          256'h8945D74087DF0566C40E28F86597C7BB7FF441A71B29B5B7686B45BB5E9358DE,
                                          256'hB41AD4941AB0E6905E5784019F32CB76BCB1CE27D85E9F39A8D71F6BC6C4331F,
                                          256'h2D3A6A125E7E25A2DDB4EB87FFEE606643AAB25E1102CAEDE0DBA59A45BAD607,
                                          256'h7C0BCCEBF1AEC76C1CFD092F710987E9C7D342F4EB0EA5C6432EFB06ACAA1C2B,
                                          256'h11C143873A8FF98885071DA3703B3D5368BBCED44FC2BCD0F7DE9CADA07D62A0,
                                          256'h5CCD82C21B84E84C968AC070913B6CA587393B31E28E204EED2ED1E2910852A7,
                                          256'h4AC8C6A79D48CF47BA068BA3B28FD6ACD57F053DC9D6A209EDBCED3E9FD450BF,
                                          256'hC650304E05A20174855D3D7B204DAD5F86ABACD131A1AB0AD39A0D5EFE2B6917,
                                          256'h3903036E09F0002AAD920BAC614D3F926FAC80DD4F16D622CA6AF643822366F6,
                                          256'hB01EDE67023E5D2BF302DE58688F6EC9AC9752B1D8CD5F1D597298810E4E385A,
                                          256'hC51999B327F52AC3D485ACB908CA5DC92CF8C6D3C6196195963981F5A2B199F6,
                                          256'h4E3038142A30251362FF6F79F2492EB6AF36B5640044C8274C9D60F6FF5E2922,
                                          256'h466D45193D2F5A27851EB344446318DE5988ED043774CD75E45D2F854FC01282,
                                          256'hBC4DE9B41D5490CA5B75AAD8EFA311FC00B3939E49D1850713CF177D312C4497,
                                          256'h4DA0A87C3DF9CA03EE0D70EBBAFEC2256737097CCE7EAD212ADCB945D92ECF5F,
                                          256'hC1423E95356CBBBA813CB486852D33E07B97D436DF617BEA021388C62A7DC86D,
                                          256'h61976CA3811120EB1FF58418D255E4446BFB5B30B1E63632F2DC624C3DCE0D0D,
                                          256'hA4E6BEFB3FE24579AA3B154991C4588CC6AA749195AB6F9DA044021089C0EA5B,
                                          256'h389D88FF194D8822E79626DE3C470409BF30523AAB56B60FBECFE33986FD3ECC,
                                          256'hCCB23289688711CA1AFCE7A6B5D2AEDC4AD0AC20372F6F2DD29EBBEBB71F5A09,
                                          256'h31254986E83195617DAD2CF9030B976FDA73F6E3CB2083586ED4629144561979,
                                          256'hDD2321A1836241052E25F6608F839236C6E6A76B952EB5716B8ACB63D66A1D6F,
                                          256'hCD1C2A4260BEE5E17CF725451E9FC36D798CBC08CC87C87E5EB6D221CB0CA87B,
                                          256'h0B07337907D0057DAE6811074F498EA0AD3CA01532861D6E26BDD9A8C2D8F90B,
                                          256'h0BFB0C192B7BF3AE7ED6DED61AD60993302E55200E38621CC574A16FBE4C09E3,
                                          256'hA6DF71896003EFA34D646F65E8DE978C604B95D0F3C2F4DFD153660035ABF919,
                                          256'hB92FD76310EF8DB5BE1161EE652268D56F4F6A517068153B5E847EB9946EB9EF,
                                          256'h91B196F95F05DBE034B2C917D0D1DBA9307F5239B0406284F9A9CCD7529C66F5,
                                          256'hB848AD6BC10DD17D6532BEB6EFA75A28EDD730657A9BEA4E57FE7B2551BE8E01,
                                          256'h35F524F324214C4CC2DFEAE418239B1F0367F8302990F102050340B1C075ED30,
                                          256'h5E05DED134063AD4B18F202C93327F0F99328C172DD2E09DCC626A0CAAD7C277,
                                          256'h7274AEED0D1CDBE71D0F707A13B560837CB577AF14A000FD354030FEE6E4A69D,
                                          256'hACE84A0B6AFDE5F9768833218589F1DBF220EBBF0A5C0DEC126B956C66248122,
                                          256'hEF95B5649B07C47F0D4624AB424E36049C40A3E31E41721ECE236145AD0D7CFF,
                                          256'h10EB0827AF406C9D4106B7096779DBF6DE770F29BFC8DDDED095A501A6F2C494,
                                          256'h80FCAB62D5AC6243202EAE66179811488E6C8EE7E2BC0A685BF4F521C2CD9ECC,
                                          256'h4137E3140FFF9B1CD52FE1BC58E01F1BBC86299A20E9CFB81E7D3E25A77F1779,
                                          256'h8D42203F6F5877C074C86D2B0FB66C234F303F1186AB32AB38630F66FA891917,
                                          256'h34C0614C9BB799AD2FAEEC155BF821319C5ABBCB60B7851D2E9C096969E90759,
                                          256'hB643CE4C863CD8FA179C53FE5A68AA21F024010A03BB37CD7C67E7975FFD6FE8,
                                          256'h92522DE360E8A9E5A875510A27123EF9AF7292745B661192E1C0CD1247D2C394,
                                          256'hEF5C168816D798C8224487868584AF0F9C31170420E50D8A4D960BF92E3C8F8A,
                                          256'hB264E9FEC44755DCB24A67E5EE43A2C689DD3D37844C79E59B820954FA9D4BE2,
                                          256'h74FD16F2234F9EB6FE74B1F3F5EB71E2F715D55BE8469F4AC40BB7D040B036F2,
                                          256'h0651E551D64CB847CCAB42864DD24792F2CCF496605891AA726DA8029A0EE875,
                                          256'hFD40E197BCFF2834A6163A4D29CC820D018E208B17B548969EBA116944FE8D3F,
                                          256'hD2A626EDDD452C3EEE676EDA0D9A387174FA00EADA48A5004BC9291ED984987C,
                                          256'h91F26300183C0BE90BF851D00142CF3FBE047BD12F6893C1C4133736BBE5B3B2,
                                          256'hF63BFDBBF4452EA520D8391BA003A6FCA9133EC40206B735B1C9867FFBFB0415,
                                          256'hBD3797F6A6F922602127825BA84473394BB7808BBE58C5F93FC181267FF6CE0E,
                                          256'hA01789F621FE5305DC59FA668BE3662A73CCABD3F850C3E3308A50B651B504D6,
                                          256'h77AF54395B0141776ADC0661BD32C972B899364A871D31318AB6C72421BCF8C6,
                                          256'h81FC858CE2A3C524F1A7218F318A20C03294496A3E28B207EB5626613345A44C,
                                          256'hFA4504FB3D05F0E2A2307BF47876E0A72291201D8533959EEA8D17F820312782,
                                          256'h0359B10D206FE69B892722071D55F08A5F7B73D7F5F77F6E641B7E688B81B867,
                                          256'h23F2F89D7D364CBABEA79F83A50254F2786104898E048A2398B4A7C114B6A234,
                                          256'h082F86AB38DD16BE2DD590E26602AFB476EBBF2040CAA73AF341C1D26BD78A51,
                                          256'h116BC61A3B38EA100E836145A48BE1DDEA75CFCFF68CDB94AEF6F8108FC328A4,
                                          256'h54D5AC7149825DB6304FE3998ED8BBB1903DB1094EC8B71132F48A87D7A91600,
                                          256'h39E79644B62F815300BBDD349EE73F04783F5C6A8E77DC2E42C50DD09B742723,
                                          256'h06A603D4087E77C5D0A10E8A50AAE92657B2BD2F40D5524E9D5088FD968799F5,
                                          256'hB73F68DB80D1C746936B4D564A665B7FF35CA3A580486EA5EE39A5E8F5B835F9,
                                          256'h6057BAD4941004DDFEC6CA3ABBCC4E3EDBA76B275A31AE86F38F29E86024086B,
                                          256'hBF9212AFEE621122E9289ADDC613B72A3556E29C43E48C716F25193DE5480AE4,
                                          256'h4002051EBB13B124CF5D034B3D03C84F9EF4EE6176FC9BFA7062FCDEC41A1766,
                                          256'h976C180E1D0D30ECC396DC414FC07179354EDCE42201796717F5A03FDF9A8834,
                                          256'hE93D307F9EF73BF5DBCA7A9E03619CB1732B90FA635BE059897963984ED61A7F,
                                          256'h5DB4EDBB34D00AD17CDB1D55F7BACF5466A89DD3C03944B982552645F8FA0184,
                                          256'h346D0A19BA19BF62E691FB960FD31642A07BAD797A099A1074AD2D0135601D2A,
                                          256'h5F50A32ADEAE4DC3CBFC26D0191C0D0C12D8638E70FDF4433C76338541CFBFC0,
                                          256'h09905A0D61DEFF51DACCE8EB2C8AB859ADF838B366B6392BB272EEA042E7900E,
                                          256'hB7EDAA849CDB4C73F0A802A65E371B5C88766C5D7D7B589C07B7E53180745D50,
                                          256'hF74A3EC14E10A49C5F30777B2CB5372C24A9AFEEB9E4D6C916E06B583F438FF6,
                                          256'h0DE432EBA133D6FA342CC161977F9CC4AD0B7CE39CD268E400C67A0D649188B5,
                                          256'h79014F7D78F974CB06E8149542EF61E072F105CD89D86D46C58CE0AE525BC193,
                                          256'h1169AE74B30BCEF2F5B295BA20CF61A730F38D84A5D23D5D08829C06D8AE19E0,
                                          256'h2385B21E9BA31773B04092B59B44CD3B5B3B27AC8186FA159004E49A53FF9EEC,
                                          256'hF63022222B89987987E75E56A4A48E3BC28CB74C0FEAF77EF6BE1725D07F743D,
                                          256'h914813055F289501615A62A60DB3AB006DD77FEC896D79F6F12AFA7555C54260,
                                          256'h8858C2003764965FBC015AC62C3A0751E5FEB9F9343EA8E623DBF205408A35B4,
                                          256'h06ADF484700072E965F4F8C2267FF81E50DB707A61A4152ACB5A780F483B04D6,
                                          256'hB6359A50EB8702ED2412CDCF6A87A9031A5D57A9F39BD37AC1095865B0BBDED9,
                                          256'hBA833077ADA35A8A9163AF64D5081F494E7D9CC2D35772FC3B726B946C246064,
                                          256'hBAAC422C46DFB676BB7555F8F8A492C6EB9CF07749DED701A15DA9A2ED5BDE1E,
                                          256'hDE4AE6948BC198D19FE8EFBDC06BA4448DBC744118FCBAE6F658DE8BB3A712D3,
                                          256'hB37081B565AE84BFC841865A8F7303446B6B76B9E253029B55A17D90DF2454DB,
                                          256'hFF3E8BB84914395195BB6CFC6E06686B3FC40E625184FB5A31320353756D80BB,
                                          256'hA9CEFE58175A8780AE838B553D5B83C2CF686EE20F7A1B8AA33673DF84181AD9,
                                          256'h8C32B70F77F5B3B385B1843640560F9851CC8AF4A1A33F80833FD53DB1DA3447,
                                          256'hEF4B04D49AD559CE73B65F21D042E7BF93CC2818E215EFE9C80DC5C3F9A24665,
                                          256'h4097D515E429EA4C48F12E7356DABDF5AF8F9D904DB3472B30D91F561FF53FDF,
                                          256'h16CBF947A22EEDB075D687C53FA9085640C3BABBB0875E9FF78691BEF14C54C8,
                                          256'hAF0DA346AAB7F5C4B14751B83DB19418A9E73DCB3FB94B95CC253AF3398B4935,
                                          256'h06D0BCB99C04A74CD1EDE4F1B783C4F56DF57504C6E0CCCAD057E8EC20203A5B,
                                          256'hAA2282207A0068EDA4E532BE5ECE57345C59B90A517E7C6833544A77CC6663C6,
                                          256'h92735E3E740042359928297D69AF61A8602C2EE23B42CC861C6A0AC9FD4E3BA2,
                                          256'h81FA45A5671FE49F4110DFA4256417A4651711CA9D0F185D8EDD7750EE6D9462,
                                          256'h3307143FBCA725305F0515C1D69DB0912E5BDF4410716B86A5872794D9569B8D,
                                          256'h450688AD8223CC7E47E6A9223106C9F21059A6B64B2363808979AD45CB4345C6,
                                          256'h58AE2FCA52D116AB733504DE198487555CA23A3D32AB7488E678719D6A83ED85,
                                          256'h041A4A60534A51CA21580035E9890660216738FDFD8D1D1164DE133F3442D39A,
                                          256'hEC20D2E5C662DD7C6E953E4249C77137ABDA61687B7871E5AC2C9AC2FE2C04B6};

   genvar                     i,j;

   generate
      for (i = 0; i < ROM_BLOCKS; i = i+1) begin : u_rom_blocks
         wire clke;

         assign clke = (i == block_addr) ? sel_i : 1'b0;

         for (j = 0; j < ROM_WORDS; j = j+1) begin : u_rom_words
            SB_RAM256x16 #(.INIT_0(ROM_DATA[256*((ROM_WORDS*(0+16*i)+j)%(16*16)) +:256]),
                           .INIT_1(ROM_DATA[256*((ROM_WORDS*(1+16*i)+j)%(16*16)) +:256]),
                           .INIT_2(ROM_DATA[256*((ROM_WORDS*(2+16*i)+j)%(16*16)) +:256]),
                           .INIT_3(ROM_DATA[256*((ROM_WORDS*(3+16*i)+j)%(16*16)) +:256]),
                           .INIT_4(ROM_DATA[256*((ROM_WORDS*(4+16*i)+j)%(16*16)) +:256]),
                           .INIT_5(ROM_DATA[256*((ROM_WORDS*(5+16*i)+j)%(16*16)) +:256]),
                           .INIT_6(ROM_DATA[256*((ROM_WORDS*(6+16*i)+j)%(16*16)) +:256]),
                           .INIT_7(ROM_DATA[256*((ROM_WORDS*(7+16*i)+j)%(16*16)) +:256]),
                           .INIT_8(ROM_DATA[256*((ROM_WORDS*(8+16*i)+j)%(16*16)) +:256]),
                           .INIT_9(ROM_DATA[256*((ROM_WORDS*(9+16*i)+j)%(16*16)) +:256]),
                           .INIT_A(ROM_DATA[256*((ROM_WORDS*(10+16*i)+j)%(16*16)) +:256]),
                           .INIT_B(ROM_DATA[256*((ROM_WORDS*(11+16*i)+j)%(16*16)) +:256]),
                           .INIT_C(ROM_DATA[256*((ROM_WORDS*(12+16*i)+j)%(16*16)) +:256]),
                           .INIT_D(ROM_DATA[256*((ROM_WORDS*(13+16*i)+j)%(16*16)) +:256]),
                           .INIT_E(ROM_DATA[256*((ROM_WORDS*(14+16*i)+j)%(16*16)) +:256]),
                           .INIT_F(ROM_DATA[256*((ROM_WORDS*(15+16*i)+j)%(16*16)) +:256]))
            u_ram256x16 (.RDATA(rdata[16*(ROM_WORDS*i+j) +:16]),
                         .RADDR(addr),
                         .RCLK(clk_i),
                         .RCLKE(clke),
                         .RE(read_i),
                         .WADDR(8'd0),
                         .WCLK(1'b0),
                         .WCLKE(1'b0),
                         .WDATA(16'b0),
                         .WE(1'b0),
                         .MASK(16'b0));
         end
      end
   endgenerate
endmodule
